module motrack

pub struct Coo {
pub mut:
	x f32
	y f32
}

pub fn track_ball(image []u8, width int, height int, nb_channels int) Coo {
	return Coo{100.0, 100.0}
}
