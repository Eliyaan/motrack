module motrack

pub struct Coord {
pub mut:
	x f32
	y f32
}

pub fn track_ball(image []u8, width int, height int, nb_channels int) Coo {
	return Coord{100.0, 100.0}
}
